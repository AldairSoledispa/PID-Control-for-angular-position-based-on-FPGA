-- SISTEMA.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SISTEMA is
	port (
		clk_clk                     : in    std_logic                     := '0';             --                    clk.clk
		clk_sdram_clk               : out   std_logic;                                        --              clk_sdram.clk
		ldr_external_interface_sclk : out   std_logic;                                        -- ldr_external_interface.sclk
		ldr_external_interface_cs_n : out   std_logic;                                        --                       .cs_n
		ldr_external_interface_dout : in    std_logic                     := '0';             --                       .dout
		ldr_external_interface_din  : out   std_logic;                                        --                       .din
		pll_locked_export           : out   std_logic;                                        --             pll_locked.export
		reset_reset_n               : in    std_logic                     := '0';             --                  reset.reset_n
		sdram_wire_addr             : out   std_logic_vector(12 downto 0);                    --             sdram_wire.addr
		sdram_wire_ba               : out   std_logic_vector(1 downto 0);                     --                       .ba
		sdram_wire_cas_n            : out   std_logic;                                        --                       .cas_n
		sdram_wire_cke              : out   std_logic;                                        --                       .cke
		sdram_wire_cs_n             : out   std_logic;                                        --                       .cs_n
		sdram_wire_dq               : inout std_logic_vector(15 downto 0) := (others => '0'); --                       .dq
		sdram_wire_dqm              : out   std_logic_vector(1 downto 0);                     --                       .dqm
		sdram_wire_ras_n            : out   std_logic;                                        --                       .ras_n
		sdram_wire_we_n             : out   std_logic                                         --                       .we_n
	);
end entity SISTEMA;

architecture rtl of SISTEMA is
	component SISTEMA_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component SISTEMA_JTAG_UART;

	component SISTEMA_LDR is
		generic (
			board          : string  := "DE10-Standard";
			board_rev      : string  := "Autodetect";
			tsclk          : integer := 0;
			numch          : integer := 0;
			max10pllmultby : integer := 0;
			max10plldivby  : integer := 0
		);
		port (
			clock       : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			waitrequest : out std_logic;                                        -- waitrequest
			read        : in  std_logic                     := 'X';             -- read
			adc_sclk    : out std_logic;                                        -- export
			adc_cs_n    : out std_logic;                                        -- export
			adc_dout    : in  std_logic                     := 'X';             -- export
			adc_din     : out std_logic                                         -- export
		);
	end component SISTEMA_LDR;

	component SISTEMA_PLL is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component SISTEMA_PLL;

	component SISTEMA_Procesador1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component SISTEMA_Procesador1;

	component SISTEMA_Procesador2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component SISTEMA_Procesador2;

	component SISTEMA_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component SISTEMA_SDRAM;

	component SISTEMA_SRAM1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component SISTEMA_SRAM1;

	component SISTEMA_SRAM2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component SISTEMA_SRAM2;

	component SISTEMA_TIMER is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component SISTEMA_TIMER;

	component SISTEMA_mm_interconnect_0 is
		port (
			PLL_outclk0_clk                               : in  std_logic                     := 'X';             -- clk
			Procesador1_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Procesador1_data_master_address               : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			Procesador1_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			Procesador1_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Procesador1_data_master_read                  : in  std_logic                     := 'X';             -- read
			Procesador1_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			Procesador1_data_master_write                 : in  std_logic                     := 'X';             -- write
			Procesador1_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Procesador1_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			Procesador1_instruction_master_address        : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			Procesador1_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			Procesador1_instruction_master_read           : in  std_logic                     := 'X';             -- read
			Procesador1_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			Procesador2_data_master_address               : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			Procesador2_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			Procesador2_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Procesador2_data_master_read                  : in  std_logic                     := 'X';             -- read
			Procesador2_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			Procesador2_data_master_write                 : in  std_logic                     := 'X';             -- write
			Procesador2_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Procesador2_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			Procesador2_instruction_master_address        : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			Procesador2_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			Procesador2_instruction_master_read           : in  std_logic                     := 'X';             -- read
			Procesador2_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			JTAG_UART_avalon_jtag_slave_address           : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write             : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read              : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect        : out std_logic;                                        -- chipselect
			LDR_adc_slave_address                         : out std_logic_vector(2 downto 0);                     -- address
			LDR_adc_slave_write                           : out std_logic;                                        -- write
			LDR_adc_slave_read                            : out std_logic;                                        -- read
			LDR_adc_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LDR_adc_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			LDR_adc_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			Procesador1_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			Procesador1_debug_mem_slave_write             : out std_logic;                                        -- write
			Procesador1_debug_mem_slave_read              : out std_logic;                                        -- read
			Procesador1_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Procesador1_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			Procesador1_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			Procesador1_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			Procesador1_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			Procesador2_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			Procesador2_debug_mem_slave_write             : out std_logic;                                        -- write
			Procesador2_debug_mem_slave_read              : out std_logic;                                        -- read
			Procesador2_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Procesador2_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			Procesador2_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			Procesador2_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			Procesador2_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			SDRAM_s1_address                              : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_s1_write                                : out std_logic;                                        -- write
			SDRAM_s1_read                                 : out std_logic;                                        -- read
			SDRAM_s1_readdata                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                            : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_s1_byteenable                           : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                        : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                           : out std_logic;                                        -- chipselect
			SRAM1_s1_address                              : out std_logic_vector(14 downto 0);                    -- address
			SRAM1_s1_write                                : out std_logic;                                        -- write
			SRAM1_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SRAM1_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			SRAM1_s1_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			SRAM1_s1_chipselect                           : out std_logic;                                        -- chipselect
			SRAM1_s1_clken                                : out std_logic;                                        -- clken
			SRAM2_s1_address                              : out std_logic_vector(14 downto 0);                    -- address
			SRAM2_s1_write                                : out std_logic;                                        -- write
			SRAM2_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SRAM2_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			SRAM2_s1_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			SRAM2_s1_chipselect                           : out std_logic;                                        -- chipselect
			SRAM2_s1_clken                                : out std_logic;                                        -- clken
			TIMER_s1_address                              : out std_logic_vector(2 downto 0);                     -- address
			TIMER_s1_write                                : out std_logic;                                        -- write
			TIMER_s1_readdata                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			TIMER_s1_writedata                            : out std_logic_vector(15 downto 0);                    -- writedata
			TIMER_s1_chipselect                           : out std_logic                                         -- chipselect
		);
	end component SISTEMA_mm_interconnect_0;

	component SISTEMA_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component SISTEMA_irq_mapper;

	component sistema_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component sistema_rst_controller;

	component sistema_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component sistema_rst_controller_001;

	signal pll_outclk0_clk                                               : std_logic;                     -- PLL:outclk_0 -> [JTAG_UART:clk, LDR:clock, Procesador1:clk, Procesador2:clk, SDRAM:clk, SRAM1:clk, SRAM2:clk, TIMER:clk, irq_mapper:clk, irq_mapper_001:clk, mm_interconnect_0:PLL_outclk0_clk, rst_controller:clk]
	signal procesador1_data_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:Procesador1_data_master_readdata -> Procesador1:d_readdata
	signal procesador1_data_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:Procesador1_data_master_waitrequest -> Procesador1:d_waitrequest
	signal procesador1_data_master_debugaccess                           : std_logic;                     -- Procesador1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Procesador1_data_master_debugaccess
	signal procesador1_data_master_address                               : std_logic_vector(26 downto 0); -- Procesador1:d_address -> mm_interconnect_0:Procesador1_data_master_address
	signal procesador1_data_master_byteenable                            : std_logic_vector(3 downto 0);  -- Procesador1:d_byteenable -> mm_interconnect_0:Procesador1_data_master_byteenable
	signal procesador1_data_master_read                                  : std_logic;                     -- Procesador1:d_read -> mm_interconnect_0:Procesador1_data_master_read
	signal procesador1_data_master_write                                 : std_logic;                     -- Procesador1:d_write -> mm_interconnect_0:Procesador1_data_master_write
	signal procesador1_data_master_writedata                             : std_logic_vector(31 downto 0); -- Procesador1:d_writedata -> mm_interconnect_0:Procesador1_data_master_writedata
	signal procesador1_instruction_master_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Procesador1_instruction_master_readdata -> Procesador1:i_readdata
	signal procesador1_instruction_master_waitrequest                    : std_logic;                     -- mm_interconnect_0:Procesador1_instruction_master_waitrequest -> Procesador1:i_waitrequest
	signal procesador1_instruction_master_address                        : std_logic_vector(26 downto 0); -- Procesador1:i_address -> mm_interconnect_0:Procesador1_instruction_master_address
	signal procesador1_instruction_master_read                           : std_logic;                     -- Procesador1:i_read -> mm_interconnect_0:Procesador1_instruction_master_read
	signal procesador2_data_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:Procesador2_data_master_readdata -> Procesador2:d_readdata
	signal procesador2_data_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:Procesador2_data_master_waitrequest -> Procesador2:d_waitrequest
	signal procesador2_data_master_debugaccess                           : std_logic;                     -- Procesador2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Procesador2_data_master_debugaccess
	signal procesador2_data_master_address                               : std_logic_vector(26 downto 0); -- Procesador2:d_address -> mm_interconnect_0:Procesador2_data_master_address
	signal procesador2_data_master_byteenable                            : std_logic_vector(3 downto 0);  -- Procesador2:d_byteenable -> mm_interconnect_0:Procesador2_data_master_byteenable
	signal procesador2_data_master_read                                  : std_logic;                     -- Procesador2:d_read -> mm_interconnect_0:Procesador2_data_master_read
	signal procesador2_data_master_write                                 : std_logic;                     -- Procesador2:d_write -> mm_interconnect_0:Procesador2_data_master_write
	signal procesador2_data_master_writedata                             : std_logic_vector(31 downto 0); -- Procesador2:d_writedata -> mm_interconnect_0:Procesador2_data_master_writedata
	signal procesador2_instruction_master_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Procesador2_instruction_master_readdata -> Procesador2:i_readdata
	signal procesador2_instruction_master_waitrequest                    : std_logic;                     -- mm_interconnect_0:Procesador2_instruction_master_waitrequest -> Procesador2:i_waitrequest
	signal procesador2_instruction_master_address                        : std_logic_vector(26 downto 0); -- Procesador2:i_address -> mm_interconnect_0:Procesador2_instruction_master_address
	signal procesador2_instruction_master_read                           : std_logic;                     -- Procesador2:i_read -> mm_interconnect_0:Procesador2_instruction_master_read
	signal mm_interconnect_0_ldr_adc_slave_readdata                      : std_logic_vector(31 downto 0); -- LDR:readdata -> mm_interconnect_0:LDR_adc_slave_readdata
	signal mm_interconnect_0_ldr_adc_slave_waitrequest                   : std_logic;                     -- LDR:waitrequest -> mm_interconnect_0:LDR_adc_slave_waitrequest
	signal mm_interconnect_0_ldr_adc_slave_address                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:LDR_adc_slave_address -> LDR:address
	signal mm_interconnect_0_ldr_adc_slave_read                          : std_logic;                     -- mm_interconnect_0:LDR_adc_slave_read -> LDR:read
	signal mm_interconnect_0_ldr_adc_slave_write                         : std_logic;                     -- mm_interconnect_0:LDR_adc_slave_write -> LDR:write
	signal mm_interconnect_0_ldr_adc_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:LDR_adc_slave_writedata -> LDR:writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_procesador1_debug_mem_slave_readdata        : std_logic_vector(31 downto 0); -- Procesador1:debug_mem_slave_readdata -> mm_interconnect_0:Procesador1_debug_mem_slave_readdata
	signal mm_interconnect_0_procesador1_debug_mem_slave_waitrequest     : std_logic;                     -- Procesador1:debug_mem_slave_waitrequest -> mm_interconnect_0:Procesador1_debug_mem_slave_waitrequest
	signal mm_interconnect_0_procesador1_debug_mem_slave_debugaccess     : std_logic;                     -- mm_interconnect_0:Procesador1_debug_mem_slave_debugaccess -> Procesador1:debug_mem_slave_debugaccess
	signal mm_interconnect_0_procesador1_debug_mem_slave_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Procesador1_debug_mem_slave_address -> Procesador1:debug_mem_slave_address
	signal mm_interconnect_0_procesador1_debug_mem_slave_read            : std_logic;                     -- mm_interconnect_0:Procesador1_debug_mem_slave_read -> Procesador1:debug_mem_slave_read
	signal mm_interconnect_0_procesador1_debug_mem_slave_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Procesador1_debug_mem_slave_byteenable -> Procesador1:debug_mem_slave_byteenable
	signal mm_interconnect_0_procesador1_debug_mem_slave_write           : std_logic;                     -- mm_interconnect_0:Procesador1_debug_mem_slave_write -> Procesador1:debug_mem_slave_write
	signal mm_interconnect_0_procesador1_debug_mem_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Procesador1_debug_mem_slave_writedata -> Procesador1:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	signal mm_interconnect_0_timer_s1_readdata                           : std_logic_vector(15 downto 0); -- TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	signal mm_interconnect_0_timer_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TIMER_s1_address -> TIMER:address
	signal mm_interconnect_0_timer_s1_write                              : std_logic;                     -- mm_interconnect_0:TIMER_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                           : std_logic_vector(15 downto 0); -- SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                        : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                            : std_logic_vector(24 downto 0); -- mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_0_sdram_s1_read                               : std_logic;                     -- mm_interconnect_0:SDRAM_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                      : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                              : std_logic;                     -- mm_interconnect_0:SDRAM_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	signal mm_interconnect_0_sram1_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:SRAM1_s1_chipselect -> SRAM1:chipselect
	signal mm_interconnect_0_sram1_s1_readdata                           : std_logic_vector(31 downto 0); -- SRAM1:readdata -> mm_interconnect_0:SRAM1_s1_readdata
	signal mm_interconnect_0_sram1_s1_address                            : std_logic_vector(14 downto 0); -- mm_interconnect_0:SRAM1_s1_address -> SRAM1:address
	signal mm_interconnect_0_sram1_s1_byteenable                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SRAM1_s1_byteenable -> SRAM1:byteenable
	signal mm_interconnect_0_sram1_s1_write                              : std_logic;                     -- mm_interconnect_0:SRAM1_s1_write -> SRAM1:write
	signal mm_interconnect_0_sram1_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:SRAM1_s1_writedata -> SRAM1:writedata
	signal mm_interconnect_0_sram1_s1_clken                              : std_logic;                     -- mm_interconnect_0:SRAM1_s1_clken -> SRAM1:clken
	signal mm_interconnect_0_procesador2_debug_mem_slave_readdata        : std_logic_vector(31 downto 0); -- Procesador2:debug_mem_slave_readdata -> mm_interconnect_0:Procesador2_debug_mem_slave_readdata
	signal mm_interconnect_0_procesador2_debug_mem_slave_waitrequest     : std_logic;                     -- Procesador2:debug_mem_slave_waitrequest -> mm_interconnect_0:Procesador2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_procesador2_debug_mem_slave_debugaccess     : std_logic;                     -- mm_interconnect_0:Procesador2_debug_mem_slave_debugaccess -> Procesador2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_procesador2_debug_mem_slave_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Procesador2_debug_mem_slave_address -> Procesador2:debug_mem_slave_address
	signal mm_interconnect_0_procesador2_debug_mem_slave_read            : std_logic;                     -- mm_interconnect_0:Procesador2_debug_mem_slave_read -> Procesador2:debug_mem_slave_read
	signal mm_interconnect_0_procesador2_debug_mem_slave_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Procesador2_debug_mem_slave_byteenable -> Procesador2:debug_mem_slave_byteenable
	signal mm_interconnect_0_procesador2_debug_mem_slave_write           : std_logic;                     -- mm_interconnect_0:Procesador2_debug_mem_slave_write -> Procesador2:debug_mem_slave_write
	signal mm_interconnect_0_procesador2_debug_mem_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Procesador2_debug_mem_slave_writedata -> Procesador2:debug_mem_slave_writedata
	signal mm_interconnect_0_sram2_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:SRAM2_s1_chipselect -> SRAM2:chipselect
	signal mm_interconnect_0_sram2_s1_readdata                           : std_logic_vector(31 downto 0); -- SRAM2:readdata -> mm_interconnect_0:SRAM2_s1_readdata
	signal mm_interconnect_0_sram2_s1_address                            : std_logic_vector(14 downto 0); -- mm_interconnect_0:SRAM2_s1_address -> SRAM2:address
	signal mm_interconnect_0_sram2_s1_byteenable                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SRAM2_s1_byteenable -> SRAM2:byteenable
	signal mm_interconnect_0_sram2_s1_write                              : std_logic;                     -- mm_interconnect_0:SRAM2_s1_write -> SRAM2:write
	signal mm_interconnect_0_sram2_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:SRAM2_s1_writedata -> SRAM2:writedata
	signal mm_interconnect_0_sram2_s1_clken                              : std_logic;                     -- mm_interconnect_0:SRAM2_s1_clken -> SRAM2:clken
	signal procesador1_irq_irq                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> Procesador1:irq
	signal procesador2_irq_irq                                           : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> Procesador2:irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- JTAG_UART:av_irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- TIMER:irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [LDR:reset, SRAM1:reset, SRAM2:reset, irq_mapper:reset, irq_mapper_001:reset, mm_interconnect_0:Procesador1_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [Procesador1:reset_req, Procesador2:reset_req, SRAM1:reset_req, SRAM2:reset_req, rst_translator:reset_req_in]
	signal procesador1_debug_reset_request_reset                         : std_logic;                     -- Procesador1:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal procesador2_debug_reset_request_reset                         : std_logic;                     -- Procesador2:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> PLL:rst
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> TIMER:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv               : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [JTAG_UART:rst_n, Procesador1:reset_n, Procesador2:reset_n, SDRAM:reset_n, TIMER:reset_n]

begin

	jtag_uart : component SISTEMA_JTAG_UART
		port map (
			clk            => pll_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	ldr : component SISTEMA_LDR
		generic map (
			board          => "DE1-SoC",
			board_rev      => "Autodetect",
			tsclk          => 8,
			numch          => 3,
			max10pllmultby => 1,
			max10plldivby  => 1
		)
		port map (
			clock       => pll_outclk0_clk,                             --                clk.clk
			reset       => rst_controller_reset_out_reset,              --              reset.reset
			write       => mm_interconnect_0_ldr_adc_slave_write,       --          adc_slave.write
			readdata    => mm_interconnect_0_ldr_adc_slave_readdata,    --                   .readdata
			writedata   => mm_interconnect_0_ldr_adc_slave_writedata,   --                   .writedata
			address     => mm_interconnect_0_ldr_adc_slave_address,     --                   .address
			waitrequest => mm_interconnect_0_ldr_adc_slave_waitrequest, --                   .waitrequest
			read        => mm_interconnect_0_ldr_adc_slave_read,        --                   .read
			adc_sclk    => ldr_external_interface_sclk,                 -- external_interface.export
			adc_cs_n    => ldr_external_interface_cs_n,                 --                   .export
			adc_dout    => ldr_external_interface_dout,                 --                   .export
			adc_din     => ldr_external_interface_din                   --                   .export
		);

	pll : component SISTEMA_PLL
		port map (
			refclk   => clk_clk,                            --  refclk.clk
			rst      => rst_controller_001_reset_out_reset, --   reset.reset
			outclk_0 => pll_outclk0_clk,                    -- outclk0.clk
			outclk_1 => clk_sdram_clk,                      -- outclk1.clk
			locked   => pll_locked_export                   --  locked.export
		);

	procesador1 : component SISTEMA_Procesador1
		port map (
			clk                                 => pll_outclk0_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                  --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                        --                          .reset_req
			d_address                           => procesador1_data_master_address,                           --               data_master.address
			d_byteenable                        => procesador1_data_master_byteenable,                        --                          .byteenable
			d_read                              => procesador1_data_master_read,                              --                          .read
			d_readdata                          => procesador1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => procesador1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => procesador1_data_master_write,                             --                          .write
			d_writedata                         => procesador1_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => procesador1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => procesador1_instruction_master_address,                    --        instruction_master.address
			i_read                              => procesador1_instruction_master_read,                       --                          .read
			i_readdata                          => procesador1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => procesador1_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => procesador1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => procesador1_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_procesador1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_procesador1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_procesador1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_procesador1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_procesador1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_procesador1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_procesador1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_procesador1_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                       -- custom_instruction_master.readra
		);

	procesador2 : component SISTEMA_Procesador2
		port map (
			clk                                 => pll_outclk0_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                  --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                        --                          .reset_req
			d_address                           => procesador2_data_master_address,                           --               data_master.address
			d_byteenable                        => procesador2_data_master_byteenable,                        --                          .byteenable
			d_read                              => procesador2_data_master_read,                              --                          .read
			d_readdata                          => procesador2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => procesador2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => procesador2_data_master_write,                             --                          .write
			d_writedata                         => procesador2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => procesador2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => procesador2_instruction_master_address,                    --        instruction_master.address
			i_read                              => procesador2_instruction_master_read,                       --                          .read
			i_readdata                          => procesador2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => procesador2_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => procesador2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => procesador2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_procesador2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_procesador2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_procesador2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_procesador2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_procesador2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_procesador2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_procesador2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_procesador2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                       -- custom_instruction_master.readra
		);

	sdram : component SISTEMA_SDRAM
		port map (
			clk            => pll_outclk0_clk,                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	sram1 : component SISTEMA_SRAM1
		port map (
			clk        => pll_outclk0_clk,                       --   clk1.clk
			address    => mm_interconnect_0_sram1_s1_address,    --     s1.address
			clken      => mm_interconnect_0_sram1_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_sram1_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_sram1_s1_write,      --       .write
			readdata   => mm_interconnect_0_sram1_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_sram1_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_sram1_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,        -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,    --       .reset_req
			freeze     => '0'                                    -- (terminated)
		);

	sram2 : component SISTEMA_SRAM2
		port map (
			clk        => pll_outclk0_clk,                       --   clk1.clk
			address    => mm_interconnect_0_sram2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_sram2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_sram2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_sram2_s1_write,      --       .write
			readdata   => mm_interconnect_0_sram2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_sram2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_sram2_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,        -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,    --       .reset_req
			freeze     => '0'                                    -- (terminated)
		);

	timer : component SISTEMA_TIMER
		port map (
			clk        => pll_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                    --   irq.irq
		);

	mm_interconnect_0 : component SISTEMA_mm_interconnect_0
		port map (
			PLL_outclk0_clk                               => pll_outclk0_clk,                                           --                             PLL_outclk0.clk
			Procesador1_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- Procesador1_reset_reset_bridge_in_reset.reset
			Procesador1_data_master_address               => procesador1_data_master_address,                           --                 Procesador1_data_master.address
			Procesador1_data_master_waitrequest           => procesador1_data_master_waitrequest,                       --                                        .waitrequest
			Procesador1_data_master_byteenable            => procesador1_data_master_byteenable,                        --                                        .byteenable
			Procesador1_data_master_read                  => procesador1_data_master_read,                              --                                        .read
			Procesador1_data_master_readdata              => procesador1_data_master_readdata,                          --                                        .readdata
			Procesador1_data_master_write                 => procesador1_data_master_write,                             --                                        .write
			Procesador1_data_master_writedata             => procesador1_data_master_writedata,                         --                                        .writedata
			Procesador1_data_master_debugaccess           => procesador1_data_master_debugaccess,                       --                                        .debugaccess
			Procesador1_instruction_master_address        => procesador1_instruction_master_address,                    --          Procesador1_instruction_master.address
			Procesador1_instruction_master_waitrequest    => procesador1_instruction_master_waitrequest,                --                                        .waitrequest
			Procesador1_instruction_master_read           => procesador1_instruction_master_read,                       --                                        .read
			Procesador1_instruction_master_readdata       => procesador1_instruction_master_readdata,                   --                                        .readdata
			Procesador2_data_master_address               => procesador2_data_master_address,                           --                 Procesador2_data_master.address
			Procesador2_data_master_waitrequest           => procesador2_data_master_waitrequest,                       --                                        .waitrequest
			Procesador2_data_master_byteenable            => procesador2_data_master_byteenable,                        --                                        .byteenable
			Procesador2_data_master_read                  => procesador2_data_master_read,                              --                                        .read
			Procesador2_data_master_readdata              => procesador2_data_master_readdata,                          --                                        .readdata
			Procesador2_data_master_write                 => procesador2_data_master_write,                             --                                        .write
			Procesador2_data_master_writedata             => procesador2_data_master_writedata,                         --                                        .writedata
			Procesador2_data_master_debugaccess           => procesador2_data_master_debugaccess,                       --                                        .debugaccess
			Procesador2_instruction_master_address        => procesador2_instruction_master_address,                    --          Procesador2_instruction_master.address
			Procesador2_instruction_master_waitrequest    => procesador2_instruction_master_waitrequest,                --                                        .waitrequest
			Procesador2_instruction_master_read           => procesador2_instruction_master_read,                       --                                        .read
			Procesador2_instruction_master_readdata       => procesador2_instruction_master_readdata,                   --                                        .readdata
			JTAG_UART_avalon_jtag_slave_address           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --             JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                        .write
			JTAG_UART_avalon_jtag_slave_read              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                        .read
			JTAG_UART_avalon_jtag_slave_readdata          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                        .readdata
			JTAG_UART_avalon_jtag_slave_writedata         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                        .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                        .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                        .chipselect
			LDR_adc_slave_address                         => mm_interconnect_0_ldr_adc_slave_address,                   --                           LDR_adc_slave.address
			LDR_adc_slave_write                           => mm_interconnect_0_ldr_adc_slave_write,                     --                                        .write
			LDR_adc_slave_read                            => mm_interconnect_0_ldr_adc_slave_read,                      --                                        .read
			LDR_adc_slave_readdata                        => mm_interconnect_0_ldr_adc_slave_readdata,                  --                                        .readdata
			LDR_adc_slave_writedata                       => mm_interconnect_0_ldr_adc_slave_writedata,                 --                                        .writedata
			LDR_adc_slave_waitrequest                     => mm_interconnect_0_ldr_adc_slave_waitrequest,               --                                        .waitrequest
			Procesador1_debug_mem_slave_address           => mm_interconnect_0_procesador1_debug_mem_slave_address,     --             Procesador1_debug_mem_slave.address
			Procesador1_debug_mem_slave_write             => mm_interconnect_0_procesador1_debug_mem_slave_write,       --                                        .write
			Procesador1_debug_mem_slave_read              => mm_interconnect_0_procesador1_debug_mem_slave_read,        --                                        .read
			Procesador1_debug_mem_slave_readdata          => mm_interconnect_0_procesador1_debug_mem_slave_readdata,    --                                        .readdata
			Procesador1_debug_mem_slave_writedata         => mm_interconnect_0_procesador1_debug_mem_slave_writedata,   --                                        .writedata
			Procesador1_debug_mem_slave_byteenable        => mm_interconnect_0_procesador1_debug_mem_slave_byteenable,  --                                        .byteenable
			Procesador1_debug_mem_slave_waitrequest       => mm_interconnect_0_procesador1_debug_mem_slave_waitrequest, --                                        .waitrequest
			Procesador1_debug_mem_slave_debugaccess       => mm_interconnect_0_procesador1_debug_mem_slave_debugaccess, --                                        .debugaccess
			Procesador2_debug_mem_slave_address           => mm_interconnect_0_procesador2_debug_mem_slave_address,     --             Procesador2_debug_mem_slave.address
			Procesador2_debug_mem_slave_write             => mm_interconnect_0_procesador2_debug_mem_slave_write,       --                                        .write
			Procesador2_debug_mem_slave_read              => mm_interconnect_0_procesador2_debug_mem_slave_read,        --                                        .read
			Procesador2_debug_mem_slave_readdata          => mm_interconnect_0_procesador2_debug_mem_slave_readdata,    --                                        .readdata
			Procesador2_debug_mem_slave_writedata         => mm_interconnect_0_procesador2_debug_mem_slave_writedata,   --                                        .writedata
			Procesador2_debug_mem_slave_byteenable        => mm_interconnect_0_procesador2_debug_mem_slave_byteenable,  --                                        .byteenable
			Procesador2_debug_mem_slave_waitrequest       => mm_interconnect_0_procesador2_debug_mem_slave_waitrequest, --                                        .waitrequest
			Procesador2_debug_mem_slave_debugaccess       => mm_interconnect_0_procesador2_debug_mem_slave_debugaccess, --                                        .debugaccess
			SDRAM_s1_address                              => mm_interconnect_0_sdram_s1_address,                        --                                SDRAM_s1.address
			SDRAM_s1_write                                => mm_interconnect_0_sdram_s1_write,                          --                                        .write
			SDRAM_s1_read                                 => mm_interconnect_0_sdram_s1_read,                           --                                        .read
			SDRAM_s1_readdata                             => mm_interconnect_0_sdram_s1_readdata,                       --                                        .readdata
			SDRAM_s1_writedata                            => mm_interconnect_0_sdram_s1_writedata,                      --                                        .writedata
			SDRAM_s1_byteenable                           => mm_interconnect_0_sdram_s1_byteenable,                     --                                        .byteenable
			SDRAM_s1_readdatavalid                        => mm_interconnect_0_sdram_s1_readdatavalid,                  --                                        .readdatavalid
			SDRAM_s1_waitrequest                          => mm_interconnect_0_sdram_s1_waitrequest,                    --                                        .waitrequest
			SDRAM_s1_chipselect                           => mm_interconnect_0_sdram_s1_chipselect,                     --                                        .chipselect
			SRAM1_s1_address                              => mm_interconnect_0_sram1_s1_address,                        --                                SRAM1_s1.address
			SRAM1_s1_write                                => mm_interconnect_0_sram1_s1_write,                          --                                        .write
			SRAM1_s1_readdata                             => mm_interconnect_0_sram1_s1_readdata,                       --                                        .readdata
			SRAM1_s1_writedata                            => mm_interconnect_0_sram1_s1_writedata,                      --                                        .writedata
			SRAM1_s1_byteenable                           => mm_interconnect_0_sram1_s1_byteenable,                     --                                        .byteenable
			SRAM1_s1_chipselect                           => mm_interconnect_0_sram1_s1_chipselect,                     --                                        .chipselect
			SRAM1_s1_clken                                => mm_interconnect_0_sram1_s1_clken,                          --                                        .clken
			SRAM2_s1_address                              => mm_interconnect_0_sram2_s1_address,                        --                                SRAM2_s1.address
			SRAM2_s1_write                                => mm_interconnect_0_sram2_s1_write,                          --                                        .write
			SRAM2_s1_readdata                             => mm_interconnect_0_sram2_s1_readdata,                       --                                        .readdata
			SRAM2_s1_writedata                            => mm_interconnect_0_sram2_s1_writedata,                      --                                        .writedata
			SRAM2_s1_byteenable                           => mm_interconnect_0_sram2_s1_byteenable,                     --                                        .byteenable
			SRAM2_s1_chipselect                           => mm_interconnect_0_sram2_s1_chipselect,                     --                                        .chipselect
			SRAM2_s1_clken                                => mm_interconnect_0_sram2_s1_clken,                          --                                        .clken
			TIMER_s1_address                              => mm_interconnect_0_timer_s1_address,                        --                                TIMER_s1.address
			TIMER_s1_write                                => mm_interconnect_0_timer_s1_write,                          --                                        .write
			TIMER_s1_readdata                             => mm_interconnect_0_timer_s1_readdata,                       --                                        .readdata
			TIMER_s1_writedata                            => mm_interconnect_0_timer_s1_writedata,                      --                                        .writedata
			TIMER_s1_chipselect                           => mm_interconnect_0_timer_s1_chipselect                      --                                        .chipselect
		);

	irq_mapper : component SISTEMA_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => procesador1_irq_irq             --    sender.irq
		);

	irq_mapper_001 : component SISTEMA_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => procesador2_irq_irq             --    sender.irq
		);

	rst_controller : component sistema_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,               -- reset_in0.reset
			reset_in1      => procesador1_debug_reset_request_reset, -- reset_in1.reset
			reset_in2      => procesador2_debug_reset_request_reset, -- reset_in2.reset
			clk            => pll_outclk0_clk,                       --       clk.clk
			reset_out      => rst_controller_reset_out_reset,        -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,    --          .reset_req
			reset_req_in0  => '0',                                   -- (terminated)
			reset_req_in1  => '0',                                   -- (terminated)
			reset_req_in2  => '0',                                   -- (terminated)
			reset_in3      => '0',                                   -- (terminated)
			reset_req_in3  => '0',                                   -- (terminated)
			reset_in4      => '0',                                   -- (terminated)
			reset_req_in4  => '0',                                   -- (terminated)
			reset_in5      => '0',                                   -- (terminated)
			reset_req_in5  => '0',                                   -- (terminated)
			reset_in6      => '0',                                   -- (terminated)
			reset_req_in6  => '0',                                   -- (terminated)
			reset_in7      => '0',                                   -- (terminated)
			reset_req_in7  => '0',                                   -- (terminated)
			reset_in8      => '0',                                   -- (terminated)
			reset_req_in8  => '0',                                   -- (terminated)
			reset_in9      => '0',                                   -- (terminated)
			reset_req_in9  => '0',                                   -- (terminated)
			reset_in10     => '0',                                   -- (terminated)
			reset_req_in10 => '0',                                   -- (terminated)
			reset_in11     => '0',                                   -- (terminated)
			reset_req_in11 => '0',                                   -- (terminated)
			reset_in12     => '0',                                   -- (terminated)
			reset_req_in12 => '0',                                   -- (terminated)
			reset_in13     => '0',                                   -- (terminated)
			reset_req_in13 => '0',                                   -- (terminated)
			reset_in14     => '0',                                   -- (terminated)
			reset_req_in14 => '0',                                   -- (terminated)
			reset_in15     => '0',                                   -- (terminated)
			reset_req_in15 => '0'                                    -- (terminated)
		);

	rst_controller_001 : component sistema_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,               -- reset_in0.reset
			reset_in1      => procesador1_debug_reset_request_reset, -- reset_in1.reset
			reset_in2      => procesador2_debug_reset_request_reset, -- reset_in2.reset
			clk            => open,                                  --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,    -- reset_out.reset
			reset_req      => open,                                  -- (terminated)
			reset_req_in0  => '0',                                   -- (terminated)
			reset_req_in1  => '0',                                   -- (terminated)
			reset_req_in2  => '0',                                   -- (terminated)
			reset_in3      => '0',                                   -- (terminated)
			reset_req_in3  => '0',                                   -- (terminated)
			reset_in4      => '0',                                   -- (terminated)
			reset_req_in4  => '0',                                   -- (terminated)
			reset_in5      => '0',                                   -- (terminated)
			reset_req_in5  => '0',                                   -- (terminated)
			reset_in6      => '0',                                   -- (terminated)
			reset_req_in6  => '0',                                   -- (terminated)
			reset_in7      => '0',                                   -- (terminated)
			reset_req_in7  => '0',                                   -- (terminated)
			reset_in8      => '0',                                   -- (terminated)
			reset_req_in8  => '0',                                   -- (terminated)
			reset_in9      => '0',                                   -- (terminated)
			reset_req_in9  => '0',                                   -- (terminated)
			reset_in10     => '0',                                   -- (terminated)
			reset_req_in10 => '0',                                   -- (terminated)
			reset_in11     => '0',                                   -- (terminated)
			reset_req_in11 => '0',                                   -- (terminated)
			reset_in12     => '0',                                   -- (terminated)
			reset_req_in12 => '0',                                   -- (terminated)
			reset_in13     => '0',                                   -- (terminated)
			reset_req_in13 => '0',                                   -- (terminated)
			reset_in14     => '0',                                   -- (terminated)
			reset_req_in14 => '0',                                   -- (terminated)
			reset_in15     => '0',                                   -- (terminated)
			reset_req_in15 => '0'                                    -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of SISTEMA
